module fragment_r_type (
    ports
);
    
endmodule